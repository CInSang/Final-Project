module
logic grid;
logic grid_evolve;

assign grid = 64'h0412_6424_0034_3C28;


    endmodule